
`ifdef RTL
    `define CYCLE_TIME 7.8
`endif
`ifdef GATE
    `define CYCLE_TIME 7.8
`endif

module PATTERN(
    // output signals
    clk,
    rst_n,
    IN_VALID_1,
    IN_VALID_2,
    ALPHA_I,
    A_I,
    D_I,
    THETA_JOINT_1,
    THETA_JOINT_2,
    THETA_JOINT_3,
    THETA_JOINT_4,
    // input signals
    OUT_VALID,
    OUT_X,
    OUT_Y,
    OUT_Z
);

//================================================================ 
//   INPUT AND OUTPUT DECLARATION
//================================================================
output reg              clk, rst_n, IN_VALID_1, IN_VALID_2;
output reg signed [5:0] ALPHA_I, THETA_JOINT_1, THETA_JOINT_2, THETA_JOINT_3, THETA_JOINT_4;
output reg        [2:0] A_I, D_I;
input                   OUT_VALID;
input      signed [10:0] OUT_X, OUT_Y, OUT_Z;

//================================================================
// parameters & integer
//================================================================
real    CYCLE = `CYCLE_TIME;
integer PATNUM = 10000;
integer patcount;
integer fin, fout;
integer lat, total_latency;
integer gap, i, cntin_num, cntout_num;
integer theta_time;
integer invalid1_rising, outvalid_rising, outvalid_falling;
real    max_err;
real    ai    [0:3];
real    di    [0:3];
real    alpha [0:2];
real    theta [0:3];
real    outx, outy, outz;
real    goldenx, goldeny, goldenz;
real    err_molecular; //no_sqrt
real    err_denominator;
real    err;

//================================================================
// clock
//================================================================
initial clk = 0;
always #(CYCLE/2.0) clk = ~clk;

//================================================================
// initial
//================================================================
initial begin
    rst_n = 1'b1;
    IN_VALID_1 = 1'b0;
    IN_VALID_2 = 1'b0;
    ALPHA_I = 6'bx;
    A_I = 3'bx;
    D_I = 3'bx;
    THETA_JOINT_1 = 6'bx;
    THETA_JOINT_2 = 6'bx;
    THETA_JOINT_3 = 6'bx;
    THETA_JOINT_4 = 6'bx;

    force clk = 0;

    total_latency = 0;
    RESET_task;

    fin = $fopen("../00_TESTBED/input.txt", "r");
    fout = $fopen("../00_TESTBED/output.txt", "r");
    max_err=0;
    for(patcount=0; patcount<PATNUM; patcount=patcount+1) begin
        lat = -1;
        invalid1_rising = 0;
        outvalid_falling = 0;
        cntin_num = $fscanf(fin, "%d", theta_time);
        //------------------------INPUT1_TASK------------------------//
        gap = $urandom_range(1, 4);  //1~5 back+1
        repeat(gap) @(negedge clk);
        IN_VALID_1 = 1'b1;
        invalid1_rising = 1;
        for(i=0; i<4; i=i+1) begin
            if(OUT_VALID!==1'b0) begin
                $display("--------------------------------------------------------------------------------------------------------------------------------------------");
                $display("                                                                           FAIL!                                                            ");
                $display("                                                     Outvalid should be 0 when Invalid_1 is high at %8t                                     ",$time);
                $display("--------------------------------------------------------------------------------------------------------------------------------------------");
                repeat(2) @(negedge clk);
                $finish;
            end

            cntin_num = $fscanf(fin, "%d", A_I);
            ai[i] = A_I;
            cntin_num = $fscanf(fin, "%d", D_I);
            di[i] = D_I;
            if(i>0) begin
                cntin_num = $fscanf(fin, "%d", ALPHA_I); 
                alpha[i-1] = ALPHA_I/32.0;
            end
            else begin
                ALPHA_I = 6'bx;
            end
            @(negedge clk);
        end

        IN_VALID_1 = 1'b0;
        ALPHA_I = 6'bx;
        A_I = 3'bx;
        D_I = 3'bx;

        err_denominator = $sqrt(ai[0]*ai[0]+di[0]*di[0])+
                          $sqrt(ai[1]*ai[1]+di[1]*di[1])+
                          $sqrt(ai[2]*ai[2]+di[2]*di[2])+
                          $sqrt(ai[3]*ai[3]+di[3]*di[3]);

        //------------------------INPUT2_TASK------------------------//
        IN_VALID_2 = 1'b1;
        for(i=0; i<theta_time; i=i+1) begin
            cntin_num = $fscanf(fin, "%d", THETA_JOINT_1);
            cntin_num = $fscanf(fin, "%d", THETA_JOINT_2);
            cntin_num = $fscanf(fin, "%d", THETA_JOINT_3);
            cntin_num = $fscanf(fin, "%d", THETA_JOINT_4);
            theta[0] = THETA_JOINT_1/32.0;
            theta[1] = THETA_JOINT_2/32.0;
            theta[2] = THETA_JOINT_3/32.0;
            theta[3] = THETA_JOINT_4/32.0;
            @(negedge clk);
        end
        IN_VALID_2 = 1'b0;
        THETA_JOINT_1 = 6'bx;
        THETA_JOINT_2 = 6'bx;
        THETA_JOINT_3 = 6'bx;
        THETA_JOINT_4 = 6'bx;

        while(!outvalid_falling) @(negedge clk);
        
    end
  
    PASS_task;
    $finish;
end


//================================================================
// always
//================================================================
always @(negedge clk) begin
    if(!OUT_VALID) begin
        if((OUT_X!==11'd0)||(OUT_Y!==11'd0)||(OUT_Z!==11'd0)) begin
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            $display("                                                                    FAIL!                                                                   ");
            $display("                                                Out should be reset after Outvalid is pulled down.                                          ");
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            repeat(3) @(negedge clk);
            $finish;
        end
    end
end

always @(negedge clk) begin
    if(invalid1_rising&&!outvalid_falling) begin
        lat = lat + 1;
        if(lat == 300) begin
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            $display("                                                                         FAIL!                                                              ");
            $display("                                                       The execution latency are over 300 cycles                                            ");
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            repeat(2) @(negedge clk);
            $finish;
        end
        @(negedge clk);
    end
    else if(outvalid_falling) begin
        total_latency = total_latency + lat;
    end
end

always @(negedge clk) begin
    if(OUT_VALID) outvalid_rising = 1;
    else if(outvalid_rising&&!OUT_VALID) outvalid_rising = 0;
    else outvalid_rising = 0;
end

always @(*) begin
    if(!OUT_VALID&&outvalid_rising) outvalid_falling = 1;
    else outvalid_falling = 0;
end

always @(negedge clk) begin
    if(OUT_VALID) begin
        if((OUT_X===11'bx)||(OUT_Y===11'bx)||(OUT_Z===11'bx)) begin
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            $display("                                                                           FAIL!                                                            ");
            $display("                                                                        OUT unknown                                                         ");
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            repeat(2) @(negedge clk);
            $finish;
        end
        cntout_num = $fscanf(fout, "%f", goldenx);
        cntout_num = $fscanf(fout, "%f", goldeny);
        cntout_num = $fscanf(fout, "%f", goldenz);
        outx = OUT_X;
        outy = OUT_Y;
        outz = OUT_Z;
        outx = outx/32.0;
        outy = outy/32.0;
        outz = outz/32.0;
        
        if((goldenx<=31.96875&&goldenx>=-32)&&(goldeny<=31.96875&&goldeny>=-32)&&(goldenz<=31.96875&&goldenz>=-32))begin
            err_molecular = (goldenx-outx)*(goldenx-outx)+
                        (goldeny-outy)*(goldeny-outy)+
                        (goldenz-outz)*(goldenz-outz)+
                        err_molecular;
			if((goldenx-outx>0.125||goldeny-outy>0.125||goldenz-outz>0.125)||(goldenx-outx<-0.125||goldeny-outy<-0.125||goldenz-outz<-0.125)) begin
				$display("%f/%f, %f/%f, %f/%f",goldenx,outx, goldeny, outy, goldenz,outz);
			end	
        end
        else begin
            err_molecular=err_molecular;
        end
    end
    else if(outvalid_falling) begin
        err = $sqrt(err_molecular/theta_time)/err_denominator;
        if(err>max_err)
            max_err=err;
        if(err>=0.015) begin
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            $display("                                                                           FAIL!                                                            ");
            $display("                                                            err rate = %f is bigger than 0.015                                              ",err);
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            repeat(2) @(negedge clk);
            $finish;
        end
        else begin
            $display("\033[0;34mPASS PATTERN NO.%4d,\033[m \033[0;32m Latency: %3d\033[m,   \033[33merr:  %f\033[0m",
                    patcount , lat, err);
        end
    end
    else if(!outvalid_falling) begin
        err_molecular = 0;
    end
end

//================================================================
// task
//================================================================

//------------------------RESET_TASK------------------------//
task RESET_task; begin
    #(0.5);    rst_n = 1'b0;

    #(3.0);
    if((OUT_VALID!==1'b0)||(OUT_X!==11'd0)||(OUT_Y!==11'd0)||(OUT_Z!==11'd0)) begin
        $display("--------------------------------------------------------------------------------------------------------------------------------------------");
        $display("                                                                         FAIL!                                                              ");
        $display("                                                  Output signal should be 0 after initial RESET at %8t ,%b,%b,%b,%b                                     ",$time,OUT_VALID,OUT_X,OUT_Y,OUT_Z);
        $display("--------------------------------------------------------------------------------------------------------------------------------------------");
        $finish;
    end
    #(14);    rst_n = 1'b1;
    #(4);     release clk; 
end endtask

task PASS_task; begin
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[30m#\033[31m#\033[30m#\033[31m#\033[31m#\033[31m#\033[31m#\033[31m#\033[30m#\033[32m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[31m#\033[31m#\033[31m#\033[32m#\033[32m#\033[31m#\033[33m#\033[35m#\033[36m#\033[35m#\033[34m#\033[31m#\033[33m#\033[36m#\033[36m#\033[34m#\033[31m#\033[31m#\033[30m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[35m#\033[36m#\033[36m#\033[35m#\033[35m#\033[33m#\033[34m#\033[35m#\033[34m#\033[35m#\033[35m#\033[32m#\033[32m#\033[31m#\033[30m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[33m#\033[36m#\033[36m#\033[34m#\033[34m#\033[35m#\033[33m#\033[32m#\033[34m#\033[35m#\033[34m#\033[35m#\033[33m#\033[31m#\033[32m#\033[32m#\033[31m#\033[30m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[33m#\033[33m#\033[35m#\033[36m#\033[35m#\033[36m#\033[36m#\033[34m#\033[33m#\033[33m#\033[33m#\033[33m#\033[34m#\033[33m#\033[35m#\033[34m#\033[34m#\033[33m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[32m#\033[33m#\033[34m#\033[35m#\033[36m#\033[35m#\033[34m#\033[34m#\033[35m#\033[35m#\033[34m#\033[34m#\033[32m#\033[32m#\033[35m#\033[32m#\033[30m#\033[34m#\033[36m#\033[35m#\033[35m#\033[34m#\033[33m#\033[31m#\033[33m#\033[34m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[32m#\033[34m#\033[35m#\033[35m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[35m#\033[36m#\033[32m#\033[30m#\033[31m#\033[31m#\033[30m#\033[34m#\033[35m#\033[34m#\033[35m#\033[35m#\033[35m#\033[35m#\033[36m#\033[36m#\033[35m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[33m#\033[35m#\033[36m#\033[35m#\033[35m#\033[36m#\033[36m#\033[35m#\033[35m#\033[35m#\033[35m#\033[35m#\033[34m#\033[35m#\033[36m#\033[35m#\033[33m#\033[31m#\033[32m#\033[34m#\033[35m#\033[35m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[36m#\033[33m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[32m#\033[35m#\033[36m#\033[35m#\033[35m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[35m#\033[36m#\033[36m#\033[36m#\033[35m#\033[33m#\033[36m#\033[36m#\033[35m#\033[35m#\033[35m#\033[35m#\033[35m#\033[35m#\033[36m#\033[36m#\033[35m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[35m#\033[36m#\033[36m#\033[35m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[35m#\033[35m#\033[35m#\033[34m#\033[35m#\033[35m#\033[36m#\033[36m#\033[33m#\033[35m#\033[36m#\033[36m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[33m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[33m#\033[36m#\033[36m#\033[35m#\033[32m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m.\033[30m.\033[30m#\033[30m#\033[31m#\033[30m#\033[31m#\033[31m#\033[32m#\033[32m#\033[33m#\033[32m#\033[33m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[33m#\033[33m#\033[34m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[35m#\033[36m#\033[36m#\033[35m#\033[31m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[31m#\033[31m#\033[31m#\033[31m#\033[31m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m.\033[34m#\033[36m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[35m#\033[36m#\033[36m#\033[35m#\033[32m#\033[30m#\033[31m#\033[31m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[31m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[31m#\033[30m#\033[33m#\033[36m#\033[35m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[31m#\033[35m#\033[36m#\033[36m#\033[36m#\033[35m#\033[30m#\033[30m#\033[31m#\033[31m#\033[31m#\033[31m#\033[31m#\033[31m#\033[31m#\033[30m#\033[30m#\033[30m#\033[31m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[30m#\033[33m#\033[35m#\033[36m#\033[33m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m#\033[32m#\033[32m#\033[32m#\033[31m#\033[34m#\033[36m#\033[36m#\033[36m#\033[36m#\033[34m#\033[31m#\033[32m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[32m#\033[31m#\033[31m#\033[30m#\033[31m#\033[30m#\033[30m#\033[30m#\033[31m#\033[30m#\033[31m#\033[34m#\033[36m#\033[36m#\033[35m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[34m#\033[32m#\033[32m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[31m#\033[30m#\033[31m#\033[30m#\033[30m#\033[30m#\033[32m#\033[35m#\033[36m#\033[36m#\033[35m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[31m#\033[32m#\033[32m#\033[31m#\033[33m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[33m#\033[32m#\033[32m#\033[32m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[31m#\033[30m#\033[30m#\033[31m#\033[33m#\033[35m#\033[36m#\033[36m#\033[35m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[31m#\033[32m#\033[32m#\033[31m#\033[33m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[34m#\033[33m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[34m#\033[35m#\033[36m#\033[36m#\033[36m#\033[34m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[31m#\033[32m#\033[32m#\033[31m#\033[33m#\033[35m#\033[36m#\033[35m#\033[35m#\033[35m#\033[35m#\033[34m#\033[34m#\033[32m#\033[32m#\033[32m#\033[33m#\033[32m#\033[31m#\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[31m#\033[31m#\033[32m#\033[31m#\033[31m#\033[30m#\033[30m#\033[30m#\033[30m.\033[32m#\033[35m#\033[36m#\033[36m#\033[36m#\033[35m#\033[33m#\033[30m#\033[31m#\033[32m#\033[31m#\033[30m.\033[31m#\033[30m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[30m#\033[30m#\033[30m.\033[30m#\033[31m#\033[31m#\033[31m#\033[31m#\033[32m#\033[31m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[32m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[34m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[31m#\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[32m#\033[35m#\033[33m#\033[32m#\033[33m#\033[34m#\033[35m#\033[30m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[32m#\033[34m#\033[35m#\033[35m#\033[35m#\033[34m#\033[33m#\033[33m#\033[33m#\033[33m#\033[33m#\033[34m#\033[35m#\033[35m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[31m#\033[31m#\033[32m#\033[35m#\033[33m#\033[33m#\033[33m#\033[33m#\033[34m#\033[34m#\033[35m#\033[35m#\033[35m#\033[35m#\033[35m#\033[34m#\033[34m#\033[31m#\033[37m.\033[31m#\033[33m#\033[34m#\033[34m#\033[34m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[32m#\033[32m#\033[31m#\033[31m#\033[31m#\033[31m#\033[32m#\033[31m#\033[35m#\033[35m#\033[33m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[31m#\033[32m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[33m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[35m#\033[35m#\033[33m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[33m#\033[32m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[34m#\033[36m#\033[35m#\033[34m#\033[34m#\033[35m#\033[35m#\033[36m#\033[36m#\033[36m#\033[35m#\033[35m#\033[35m#\033[34m#\033[32m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m#\033[30m#\033[30m#\033[37m.\033[30m.\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[34m#\033[36m#\033[36m#\033[35m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[34m#\033[32m#\033[33m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[34m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m#\033[30m#\033[30m#\033[37m.\033[30m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[33m#\033[34m#\033[35m#\033[36m#\033[36m#\033[36m#\033[35m#\033[35m#\033[35m#\033[33m#\033[32m#\033[31m#\033[34m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[32m#\033[32m#\033[33m#\033[33m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[33m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[30m.\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[31m#\033[31m#\033[31m#\033[31m#\033[30m#\033[30m#\033[30m#\033[33m#\033[35m#\033[36m#\033[36m#\033[35m#\033[34m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[34m#\033[33m#\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[31m#\033[30m#\033[30m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[32m#\033[32m#\033[31m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[34m#\033[36m#\033[35m#\033[31m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[30m#\033[30m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[35m#\033[36m#\033[36m#\033[35m#\033[32m#\033[32m#\033[32m#\033[32m#\033[32m#\033[31m#\033[31m#\033[30m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[35m#\033[34m#\033[33m#\033[33m#\033[30m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[33m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[34m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[30m.\033[33m#\033[35m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[36m#\033[33m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[31m#\033[33m#\033[33m#\033[34m#\033[34m#\033[33m#\033[32m#\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.\033[37m.");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                 Congratulations!                                                     ");
    $display("                                           You have passed all patterns!                                              ");
    $display("                                           Your execution cycles = %5d cycles                                         ", total_latency);
    $display("                                           Your clock period = %.1f ns                                                ", CYCLE);
    $display("                                           Your total latency = %.1f ns                                               ", total_latency*CYCLE);
    $display("                                           Your max   error  = %.10f                                                ", max_err);
    $display("----------------------------------------------------------------------------------------------------------------------");
    $finish;
end endtask



endmodule